package pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  //`include "design.sv"
  `include "sequence_item.sv"
  `include "sequencer.sv"
  `include "sequence.sv"
  `include "driver.sv"
  `include "coverage.sv"
  `include "monitor.sv"
  `include "agent.sv"
  `include "scoreboard.sv"
  `include "environment.sv"
  `include "test.sv" 
  //`include "test_2.sv"

endpackage : pkg
