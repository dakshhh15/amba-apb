package pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"
  `include "sequence_item.sv"
  `include "reset_seq.sv"
  `include "main_seq.sv"
  `include "sequencer.sv"
  `include "coverage.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "agent.sv"
  `include "scoreboard.sv"
  `include "environment.sv"
  `include "test.sv" 

endpackage : pkg
